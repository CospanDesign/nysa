
/*
  METADATA

  DRT_ID:${DRT_ID}
  DRT_FLAGS:${DRT_FLAGS}
  DRT_SIZE:${DRT_SIZE}
*/

module ${NAME} (
);

endmodule
