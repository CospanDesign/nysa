// top.v

${LICENSE}

/*

  Description:
    Top file for a Nysa IBuilder Project.

  Author: Dave McCoy dave.mccoy@cospandesign.com

  ***WARNING***
  
  THIS FILE IS AUTOMATICALLY GENERATED! ANY CHANGES MADE DIRECTLY WILL BE
  OVERWRITTEN WHEN REGENERATED
  
*/



/*
Log:
5/19/2013:
  -Initial version of template based top file. (Previous versions were
    completely procedurally generated)
*/

module top (
${PORTS}
);

//Local Parameters
${LOCAL_PARAMS}
//Registers/Wires
${SIGNALS}
//Submodules

//Host Interface
${HOST_INTERFACE}

//Master
${MASTER}

//Peripheral Interconnect
${INTERCONNECT}

//Memory Interconnect
${MEM_INTERCONNECT}

//Peripheral Slaves
${SLAVES}

//Memory Slaves
${MEMORY_SLAVES}

//Asynchronous Logic
${ASSYNCHRONOUS_LOGIC}

//Synchronous Logic
${SYNCHRONOUS_LOGIC}


endmodule
