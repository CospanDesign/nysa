module ();

endmodule
